interface intf;
  
endinterface