package pack_mem;
    `include "transaction.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "scoreboard.sv"
    `include "subscriber.sv"
    `include "env.sv"
endpackage